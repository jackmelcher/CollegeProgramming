module rom_tb;
	reg[31:0] addr;
	wire[31:0] dataIO;
	
rom L1(
	.addr(addr)
  ,.dataIO(dataIO)
);

initial begin
	addr = 32'b00000000000000000000000000000000;
	#100;
	
	addr = 32'b00000000000000000000000000000001;
	#100;
	
	addr = 32'b00000000000000000000000000000010;
	#100;
	
	addr = 32'b00000000000000000000000000000011;
	#100;
	
	addr = 32'b00000000000000000000000000000100;
	#100;
	
	addr = 32'b00000000000000000000000000000101;
	#100;
	
end
endmodule